
module object

pub struct Object {
pub:
	vertices  []f32
	textures  []f32
	normals   []f32
}